module blind(
	input i_clk,
	input i_rst,
	input i_start,
	output oHD,
	output oVD,
	output oDEN,
	output [7:0] oR,
	output [7:0] oG,
	output [7:0] oB
);